`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.07.2025 09:35:48
// Design Name: 
// Module Name: FOMUX_Using_TOMUX_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FOMUX_Using_TOMUX_TB;
reg a,b,c,d,s0,s1;
wire out;
FOMUX_Using_TOMUX uut(a,b,c,d,s1,s0);
initial begin
s1=0;s0=0;a=1;b=0;c=0;d=0;
#10
s1=0;s0=1;a=0;b=1;c=0;d=0;
#10
s1=1;s0=0;a=1;b=0;c=1;d=0;
#10
s1=1;s0=1;a=1;b=0;c=0;d=1;
#10
$finish();
end
endmodule
