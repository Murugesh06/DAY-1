`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.07.2025 11:07:13
// Design Name: 
// Module Name: fa_using_nand
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fa_using_nand(input a,b,c,output s,ca);
wire w1,w2,w3,w4,w5,w6,w7;
nand(w1,a,b);
nand(w2,a,w1);
nand(w3,w1,b);
nand(w4,w2,w3);
nand(w5,w4,c);
nand(w6,w4,w5);
nand(w7,w5,c);
nand(s,w6,w7);
nand(ca,w7,w1);
endmodule
